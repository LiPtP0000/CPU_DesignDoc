module CAR (
    i_clk,
    i_rst_n
);
    
endmodule