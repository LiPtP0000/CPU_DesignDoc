/*
module TOP
Author: LiPtP

Should instantiate:
1. CPU
2. User Interface

This is the very top module of the CPU.
*/