/*
module CPU_TOP
Author: LiPtP

Should instantiate:
1. External Bus
2. Control Unit
3. Internal Registers
4. Memories
and they should be at the same hierarchy level as they explains the whole CPU. 

The user interface should acknowledge part of CPU status and provide input to CPU, so it should be at the same level as this module.

*/